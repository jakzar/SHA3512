library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.env.stop;

entity tb_sha3_512_iota_fun is
end tb_sha3_512_iota_fun;

architecture behavior of tb_sha3_512_iota_fun is
    signal in_data  : std_logic_vector(1599 downto 0);
    signal in_RC  : std_logic_vector(63 downto 0);
    signal out_data : std_logic_vector(1599 downto 0);
begin
    uut: entity work.sha3_512_iota_fun port map(in_data, in_RC, out_data);
    process
    begin
        --dane do przetworzenia przed przeksztalceniem iota w pierwszej rundzie dla wiadomosci o dlugosci 0 bitow zgodnie z wektorami testowymi oraz wartosc RC (LE)
        in_data <= x"0600000000080000000000000060000000200300000800000600000000000000002003000060000000000000000000000000C80000C0000000000000000000200000000000C000000000C800000000200C00000000000000C00C00000000000000000000000000008C0C00000000000040000000000000000018006400000000008000000000000000180000000000000080006400000000000000000000000000000000400600400000000000004000180000004006000000000000000000401800000000004000";
        in_RC<=x"0100000000000000";
        wait for 10 ns;
        if(out_data = x"0700000000080000000000000060000000200300000800000600000000000000002003000060000000000000000000000000C80000C0000000000000000000200000000000C000000000C800000000200C00000000000000C00C00000000000000000000000000008C0C00000000000040000000000000000018006400000000008000000000000000180000000000000080006400000000000000000000000000000000400600400000000000004000180000004006000000000000000000401800000000004000") then
            report "Iota is correct";
        else
            report "Iota is incorrect";
        end if;
        
        --dane do przetworzenia przed przeksztalceniem iota w 23 rundzie dla wiadomosci o dlugosci 0 bitow zgodnie z wektorami testowymi oraz wartosc RC (LE)
        in_data <= x"AE1F734CA23A9A45C8B567DC185A756E97C982164FE25859E0D1DCC1475C80A615B2123AF1F5F94C11E3E9402C3AC558F500199D95B6D3E301758586281DCD26364BC5B8E78F53B823DDA7F4DE9FAD00E67DB72F9F9FEA0CE3C9FEF15A76ADC585EB2EFD1187FB65F9C9A273315167E314FA68B6A322D407015D502ACDEC8C885C4F7784CED04609BB35154A96484B5625D3417C88607ACDE4C2C99BAE5EDF9EEA2AD0FB55A226189E11D24960433E2B0EE045A473099776DD5DE739DB9BA819D54CB903A7A5D7EE";
        in_RC<=x"0880008000000080";
        wait for 10 ns;
        if(out_data = x"A69F73CCA23A9AC5C8B567DC185A756E97C982164FE25859E0D1DCC1475C80A615B2123AF1F5F94C11E3E9402C3AC558F500199D95B6D3E301758586281DCD26364BC5B8E78F53B823DDA7F4DE9FAD00E67DB72F9F9FEA0CE3C9FEF15A76ADC585EB2EFD1187FB65F9C9A273315167E314FA68B6A322D407015D502ACDEC8C885C4F7784CED04609BB35154A96484B5625D3417C88607ACDE4C2C99BAE5EDF9EEA2AD0FB55A226189E11D24960433E2B0EE045A473099776DD5DE739DB9BA819D54CB903A7A5D7EE") then
            report "Iota is correct";
        else
            report "Iota is incorrect";
        end if;

        --dane do przetworzenia przed przeksztalceniem iota w pierwszej rundzi dla wiadomosci o dlugosci 1630 bitow zgodnie z wektorami testowymi oraz wartosc RC (LE)
        in_data <= x"0000000000000000D2D2D2D2D2D2D2D20000000000000000E8E8E8E8E8E8E8E83A3A3A3A3A3A3A3A535353535353535300000000000000001D1D1D1D1D1D1D1D4E4E4E4E4E4E4E4E00000000000000004141414141414141E8E8E8E8E8E8E8E80000000000000000414141414141414126262626262626261D1D1D1D1D1D1D1D0000000000000000474747474747474718181818181818184747474747474747E8E8E8E8E8E8E8E835353535353535350000000000000000AFAFAFAFAFAFAFAF1212121212121212";
        in_RC<=x"0100000000000000";
        wait for 10 ns;
        if(out_data = x"0100000000000000D2D2D2D2D2D2D2D20000000000000000E8E8E8E8E8E8E8E83A3A3A3A3A3A3A3A535353535353535300000000000000001D1D1D1D1D1D1D1D4E4E4E4E4E4E4E4E00000000000000004141414141414141E8E8E8E8E8E8E8E80000000000000000414141414141414126262626262626261D1D1D1D1D1D1D1D0000000000000000474747474747474718181818181818184747474747474747E8E8E8E8E8E8E8E835353535353535350000000000000000AFAFAFAFAFAFAFAF1212121212121212") then
            report "Iota is correct";
        else
            report "Iota is incorrect";
        end if;
        stop;
    end process;

end behavior;
