library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.env.stop;

entity tb_sha3_512_theta_fun is
end tb_sha3_512_theta_fun;

architecture behavior of tb_sha3_512_theta_fun is
    signal in_data  : std_logic_vector(1599 downto 0);
    signal out_data : std_logic_vector(1599 downto 0);

begin
    uut: entity work.sha3_512_theta_fun port map(in_data, out_data);
    process
    begin
        wait for 10 ns;
        --dane do przetworzenia przed przeksztalceniem theta w pierwszej rundzie dla wiadomosci o dlugosci 0 bitow zgodnie z wektorami testowymi
        in_data <= x"0600000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
        wait for 10 ns;
        if(out_data = x"06000000000000000600000000000000010000000000000000000000000000000C0000000000008000000000000000000600000000000000010000000000000000000000000000800C0000000000008000000000000000000600000000000000010000000000000000000000000000000C0000000000008000000000000000000600000000000000010000000000000000000000000000000C0000000000008000000000000000000600000000000000010000000000000000000000000000000C00000000000080") then
            report "Hash is correct";
        else
            report "Hash is incorrect";
        end if;
        
        --dane do przetworzenia przed przeksztalceniem theta w 23 rundzie dla wiadomosci o dlugosci 0 bitow zgodnie z wektorami testowymi
        in_data <= x"05E970FDF2F2E59C31145914C5A146AD8EE71F4FFE304EBC8DB291A1AFCAC250C4A158255AC01EF4A1D98419E2B17CB1B62D8E1F607B975A1373A7E30EADEA7A095CDE8FAA3B951939D480B43F569E9F9140758913E8D3CC0FCC10AB5B9DC3F3ACE42B48EE9933E3B16B00DA0A2B5EE3B25EA0B8C3DF5F60E1780F6A5818CD055F82B54EA07A2FC487F4DAB902139B63649E707D0EAE9098A4CBB7884E2BD894216533D18298FCD6F6F064C7C95323882D63D6B595D5B882D33E8081B1477CD900526162717644C7";
        wait for 10 ns;
        if(out_data = x"AC55F36C453B9A54F3B6DB130F0F5416AA2B777709399A23C03053CE1521F024AC5F9D8059A40D7B0865078855780379748F0C18AAD585E137BFCFDBF9A43EE544DE1CE010D0A76D512A45113C328D1038FCF618A421AC04CD6E92AC9133D148882843701990E77CFCE9C2B5B0C06C97DAA0651DC0BB4CEF48C48CFBEFD1B2CD9D2037496AD43D7FA338B281F51A4FFC291CB212B445A2ECCC35722D4D4FCB1B88D9B0403551831E3452E6C003FD313309AFBE8D62DC6C1D9EBC42EE0BAC4EAD68ACA4C772125748") then
            report "Hash is correct";
        else
            report "Hash is incorrect";
        end if;
        --dane do przetworzenia przed przeksztalceniem theta w pierwszej rundzi dla wiadomosci o dlugosci 1630 bitow zgodnie z wektorami testowymi
        in_data <= x"A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A30000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
        wait for 10 ns;
        if(out_data = x"0000000000000000A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3E4E4E4E4E4E4E4E4A3A3A3A3A3A3A3A30000000000000000A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3E4E4E4E4E4E4E4E40000000000000000A3A3A3A3A3A3A3A30000000000000000000000000000000047474747474747470000000000000000A3A3A3A3A3A3A3A30000000000000000000000000000000047474747474747470000000000000000A3A3A3A3A3A3A3A30000000000000000000000000000000047474747474747470000000000000000") then
            report "Hash is correct";
        else
            report "Hash is incorrect";
        end if;
        stop;
    end process;

end behavior;
