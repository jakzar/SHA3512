library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.env.stop;

entity tb_sha3_512_round_fun is
end tb_sha3_512_round_fun;

architecture behavior of tb_sha3_512_round_fun is
    signal in_data  : std_logic_vector(1599 downto 0);
    signal in_RC  : std_logic_vector(63 downto 0);
    signal out_data : std_logic_vector(1599 downto 0);

begin
    uut: entity work.sha3_512_round_fun port map(in_data, in_RC, out_data);
    process
    begin
        --dane do przetworzenia przed przeksztalceniem pierwszej rundy dla wiadomosci o dlugosci 0 bitow zgodnie z wektorami testowymi oraz wartosc RC (LE)
        in_data <= x"0600000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
        in_RC<=x"0100000000000000";
        wait for 10 ns;
        if(out_data = x"0700000000080000000000000060000000200300000800000600000000000000002003000060000000000000000000000000C80000C0000000000000000000200000000000C000000000C800000000200C00000000000000C00C00000000000000000000000000008C0C00000000000040000000000000000018006400000000008000000000000000180000000000000080006400000000000000000000000000000000400600400000000000004000180000004006000000000000000000401800000000004000") then
            report "Round value is correct";
        else
            report "Round value is incorrect";
        end if;
        
        --dane do przetworzenia przed przeksztalceniem w 23 rundzie dla wiadomosci o dlugosci 0 bitow zgodnie z wektorami testowymi oraz wartosc RC (LE)
        in_data <= x"05E970FDF2F2E59C31145914C5A146AD8EE71F4FFE304EBC8DB291A1AFCAC250C4A158255AC01EF4A1D98419E2B17CB1B62D8E1F607B975A1373A7E30EADEA7A095CDE8FAA3B951939D480B43F569E9F9140758913E8D3CC0FCC10AB5B9DC3F3ACE42B48EE9933E3B16B00DA0A2B5EE3B25EA0B8C3DF5F60E1780F6A5818CD055F82B54EA07A2FC487F4DAB902139B63649E707D0EAE9098A4CBB7884E2BD894216533D18298FCD6F6F064C7C95323882D63D6B595D5B882D33E8081B1477CD900526162717644C7";
        in_RC<=x"0880008000000080";
        wait for 10 ns;
        if(out_data = x"A69F73CCA23A9AC5C8B567DC185A756E97C982164FE25859E0D1DCC1475C80A615B2123AF1F5F94C11E3E9402C3AC558F500199D95B6D3E301758586281DCD26364BC5B8E78F53B823DDA7F4DE9FAD00E67DB72F9F9FEA0CE3C9FEF15A76ADC585EB2EFD1187FB65F9C9A273315167E314FA68B6A322D407015D502ACDEC8C885C4F7784CED04609BB35154A96484B5625D3417C88607ACDE4C2C99BAE5EDF9EEA2AD0FB55A226189E11D24960433E2B0EE045A473099776DD5DE739DB9BA819D54CB903A7A5D7EE") then
            report "Round value is correct";
        else
            report "Round value is incorrect";
        end if;

        --dane do przetworzenia przed przeksztalceniem pierwszej rundy dla wiadomosci o dlugosci 1630 bitow zgodnie z wektorami testowymi oraz wartosc RC (LE)
        in_data <= x"A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A30000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
        in_RC<=x"0100000000000000";
        wait for 10 ns;
        if(out_data = x"0100000000000000D2D2D2D2D2D2D2D20000000000000000E8E8E8E8E8E8E8E83A3A3A3A3A3A3A3A535353535353535300000000000000001D1D1D1D1D1D1D1D4E4E4E4E4E4E4E4E00000000000000004141414141414141E8E8E8E8E8E8E8E80000000000000000414141414141414126262626262626261D1D1D1D1D1D1D1D0000000000000000474747474747474718181818181818184747474747474747E8E8E8E8E8E8E8E835353535353535350000000000000000AFAFAFAFAFAFAFAF1212121212121212") then
            report "Round value is correct";
        else
            report "Round value is incorrect";
        end if;
        stop;
    end process;

end behavior;
