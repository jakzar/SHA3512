library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.env.stop;

entity tb_sha3_512_pi_fun is
end tb_sha3_512_pi_fun;

architecture behavior of tb_sha3_512_pi_fun is
    signal in_data  : std_logic_vector(1599 downto 0);
    signal out_data : std_logic_vector(1599 downto 0);

begin
    uut: entity work.sha3_512_pi_fun port map(in_data, out_data);
    process
    begin
        --dane do przetworzenia przed przeksztalceniem pi w pierwszej rundzie dla wiadomosci o dlugosci 0 bitow zgodnie z wektorami testowymi
        in_data <= x"06000000000000000C0000000000000000000000000000400000000000000000000000640000000000000000000000000000000000600000400000000000000000000000000040000000C800000000000000000000000000001800000000000000000000000800000000000000000000000000004006000000000000000000000000000000C0000000800000000000000000000000000000800C00000000000000000000000000001800000000000000000000000000002000000000000000000020030000000000";
        wait for 10 ns;
        if(out_data = x"0600000000000000000000000060000000000000000800000000000000000000002003000000000000000000000000000000C8000000000000000000000000000000000000C0000000000000000000200C0000000000000040000000000000000000000000000000800C00000000000000000000000000000000006400000000000000000000000000180000000000000080000000000000000000000000000000000000000000400000000000004000000000004006000000000000000000001800000000000000") then
            report "Pi is correct";
        else
            report "Pi is incorrect";
        end if;
        
        --dane do przetworzenia przed przeksztalceniem pi w 23 rundzie dla wiadomosci o dlugosci 0 bitow zgodnie z wektorami testowymi
        in_data <= x"AC55F36C453B9A54E66DB7271E1EA82CEACADD5D428EE68811024F020C33E55C226DD863FDEA04CC588537908750768080A15A5D184EF7C8F9CDEFF3763EA94F6F0E7008E8D33622D30811A55214C123C0E1B7C7200D61252335BB49B246CE4482CB803CE743441981D92EF9D3856B610EE05DA6776DD0B2F7DFA3659B91881926498DBAE7AF13E427FE511CD9C07A8D48943D85435682B61BCC35722D4D4FCB0D7A2066C302D544D04899030FF4C7CCE1D5B7518C9BAD23BC42EE0BAC4EAD9E15121A2BE9B19CC4";
        wait for 10 ns;
        if(out_data = x"AC55F36C453B9A5480A15A5D184EF7C882CB803CE743441948943D85435682B615121A2BE9B19CC411024F020C33E55CD30811A55214C123C0E1B7C7200D612526498DBAE7AF13E4E1D5B7518C9BAD23E66DB7271E1EA82CF9CDEFF3763EA94F81D92EF9D3856B611BCC35722D4D4FCB0D7A2066C302D544226DD863FDEA04CC58853790875076802335BB49B246CE4427FE511CD9C07A8DBC42EE0BAC4EAD9EEACADD5D428EE6886F0E7008E8D336220EE05DA6776DD0B2F7DFA3659B918819D04899030FF4C7CC") then
            report "Pi is correct";
        else
            report "Pi is incorrect";
        end if;
        --dane do przetworzenia przed przeksztalceniem pi w pierwszej rundzi dla wiadomosci o dlugosci 1630 bitow zgodnie z wektorami testowymi
        in_data <= x"00000000000000004747474747474747E8E8E8E8E8E8E8E84E4E4E4E4E4E4E4E1D1D1D1D1D1D1D1D00000000000000003A3A3A3A3A3A3A3AE8E8E8E8E8E8E8E8727272727272727200000000000000001D1D1D1D1D1D1D1D000000000000000000000000000000008E8E8E8E8E8E8E8E0000000000000000474747474747474700000000000000000000000000000000E8E8E8E8E8E8E8E800000000000000008E8E8E8E8E8E8E8E0000000000000000000000000000000047474747474747470000000000000000";
        wait for 10 ns;
        if(out_data = x"00000000000000003A3A3A3A3A3A3A3A0000000000000000E8E8E8E8E8E8E8E800000000000000004E4E4E4E4E4E4E4E00000000000000001D1D1D1D1D1D1D1D000000000000000000000000000000004747474747474747E8E8E8E8E8E8E8E88E8E8E8E8E8E8E8E00000000000000008E8E8E8E8E8E8E8E1D1D1D1D1D1D1D1D0000000000000000000000000000000000000000000000004747474747474747E8E8E8E8E8E8E8E87272727272727272000000000000000047474747474747470000000000000000") then
            report "Pi is correct";
        else
            report "Pi is incorrect";
        end if;
        stop;
    end process;

end behavior;
