library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.env.stop;

entity tb_sha3_512_rho_fun is
end tb_sha3_512_rho_fun;

architecture behavior of tb_sha3_512_rho_fun is
    signal in_data  : std_logic_vector(1599 downto 0);
    signal out_data : std_logic_vector(1599 downto 0);


begin
    uut: entity work.sha3_512_rho_fun port map(in_data, out_data);
    process
    begin
        --dane do przetworzenia przed przeksztalceniem rho w pierwszej rundzie dla wiadomosci o dlugosci 0 bitow zgodnie z wektorami testowymi
        in_data <= x"06000000000000000600000000000000010000000000000000000000000000000C0000000000008000000000000000000600000000000000010000000000000000000000000000800C0000000000008000000000000000000600000000000000010000000000000000000000000000000C0000000000008000000000000000000600000000000000010000000000000000000000000000000C0000000000008000000000000000000600000000000000010000000000000000000000000000000C00000000000080";
        wait for 10 ns;
        if(out_data = x"06000000000000000C0000000000000000000000000000400000000000000000000000640000000000000000000000000000000000600000400000000000000000000000000040000000C800000000000000000000000000001800000000000000000000000800000000000000000000000000004006000000000000000000000000000000C0000000800000000000000000000000000000800C00000000000000000000000000001800000000000000000000000000002000000000000000000020030000000000") then
            report "Rho is correct";
        else
            report "Rho is incorrect";
        end if;
        
        --dane do przetworzenia przed przeksztalceniem rho w 23 rundzie dla wiadomosci o dlugosci 0 bitow zgodnie z wektorami testowymi
        in_data <= x"AC55F36C453B9A54F3B6DB130F0F5416AA2B777709399A23C03053CE1521F024AC5F9D8059A40D7B0865078855780379748F0C18AAD585E137BFCFDBF9A43EE544DE1CE010D0A76D512A45113C328D1038FCF618A421AC04CD6E92AC9133D148882843701990E77CFCE9C2B5B0C06C97DAA0651DC0BB4CEF48C48CFBEFD1B2CD9D2037496AD43D7FA338B281F51A4FFC291CB212B445A2ECCC35722D4D4FCB1B88D9B0403551831E3452E6C003FD313309AFBE8D62DC6C1D9EBC42EE0BAC4EAD68ACA4C772125748";
        wait for 10 ns;
        if(out_data = x"AC55F36C453B9A54E66DB7271E1EA82CEACADD5D428EE68811024F020C33E55C226DD863FDEA04CC588537908750768080A15A5D184EF7C8F9CDEFF3763EA94F6F0E7008E8D33622D30811A55214C123C0E1B7C7200D61252335BB49B246CE4482CB803CE743441981D92EF9D3856B610EE05DA6776DD0B2F7DFA3659B91881926498DBAE7AF13E427FE511CD9C07A8D48943D85435682B61BCC35722D4D4FCB0D7A2066C302D544D04899030FF4C7CCE1D5B7518C9BAD23BC42EE0BAC4EAD9E15121A2BE9B19CC4") then
            report "Rho is correct";
        else
            report "Rho is incorrect";
        end if;
        --dane do przetworzenia przed przeksztalceniem rho w pierwszej rundzi dla wiadomosci o dlugosci 1630 bitow zgodnie z wektorami testowymi
        in_data <= x"0000000000000000A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3E4E4E4E4E4E4E4E4A3A3A3A3A3A3A3A30000000000000000A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3E4E4E4E4E4E4E4E40000000000000000A3A3A3A3A3A3A3A30000000000000000000000000000000047474747474747470000000000000000A3A3A3A3A3A3A3A30000000000000000000000000000000047474747474747470000000000000000A3A3A3A3A3A3A3A30000000000000000000000000000000047474747474747470000000000000000";
        wait for 10 ns;
        if(out_data = x"00000000000000004747474747474747E8E8E8E8E8E8E8E84E4E4E4E4E4E4E4E1D1D1D1D1D1D1D1D00000000000000003A3A3A3A3A3A3A3AE8E8E8E8E8E8E8E8727272727272727200000000000000001D1D1D1D1D1D1D1D000000000000000000000000000000008E8E8E8E8E8E8E8E0000000000000000474747474747474700000000000000000000000000000000E8E8E8E8E8E8E8E800000000000000008E8E8E8E8E8E8E8E0000000000000000000000000000000047474747474747470000000000000000") then
            report "Hash is correct";
        else
            report "Hash is incorrect";
        end if;
        stop;
    end process;

end behavior;
